module test(
input reg a, b,
output reg c);
reg tempa;
 always @(b)begin
a <= !a;
c <= b;
end
endmodule 